LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.BasicPackage.ALL;

PACKAGE ImagePackage IS

TYPE ImageMatrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_logic_vector(3 DOWNTO 0);

CONSTANT spaceshipR : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"4" , x"4" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"9" , x"9" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"6" , x"1" , x"1" , x"6" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"1" , x"2" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"2" , x"1" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"0" , x"0" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"3" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"6" , x"B" , x"B" , x"9" , x"9" , x"B" , x"B" , x"6" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"5" , x"3" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"8" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"8" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"3" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"1" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"4" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"4" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"1" , x"1" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"3" , x"3" , x"3" , x"3" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"F" , x"F" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT spaceshipG : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"5" , x"5" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"8" , x"8" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"5" , x"1" , x"1" , x"6" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"1" , x"2" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"2" , x"1" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"A" , x"A" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"3" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"6" , x"B" , x"B" , x"8" , x"8" , x"B" , x"B" , x"6" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"5" , x"3" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"8" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"8" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"3" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"1" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"4" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"4" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"3" , x"3" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"1" , x"1" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"3" , x"3" , x"3" , x"3" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"C" , x"7" , x"7" , x"C" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"C" , x"F" , x"7" , x"C" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"7" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"C" , x"C" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"C" , x"C" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT spaceshipB : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"3" , x"3" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"9" , x"9" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"6" , x"1" , x"1" , x"6" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"1" , x"1" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"1" , x"1" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"2" , x"E" , x"E" , x"2" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"4" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"4" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"6" , x"B" , x"B" , x"9" , x"9" , x"B" , x"B" , x"6" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"5" , x"4" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"8" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"8" , x"D" , x"D" , x"D" , x"D" , x"D" , x"D" , x"4" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"1" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"6" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"6" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"4" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"4" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"4" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"6" , x"3" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"4" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"4" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"3" , x"6" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"4" , x"4" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"B" , x"B" , x"1" , x"1" , x"B" , x"B" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"4" , x"4" , x"4" , x"4" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"2" , x"2" , x"0" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"0" , x"2" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT BackgroundR : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"3" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"3" , x"3" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"3" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"1" , x"3" , x"3" , x"3" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"3" , x"4" , x"3" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"3" , x"4" , x"3" , x"3" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"4" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" ),
( x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" ),
( x"1" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" ),
( x"1" , x"2" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"4" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"4" , x"3" , x"2" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"3" , x"4" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"4" , x"4" , x"3" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"3" , x"3" , x"4" , x"3" , x"4" , x"3" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"4" , x"4" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT BackgroundG : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"2" , x"3" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" ),
( x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" ),
( x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" ),
( x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT BackgroundB : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"3" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"3" , x"3" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" ),
( x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"3" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"1" , x"3" , x"3" , x"3" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" ),
( x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"3" , x"3" , x"3" , x"2" , x"2" , x"1" , x"2" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" ),
( x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" ),
( x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"1" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"1" , x"2" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"2" , x"3" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" ),
( x"2" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"2" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_5R : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"F" , x"F" , x"2" , x"F" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"A" , x"A" , x"A" , x"F" , x"F" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"F" , x"F" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"A" , x"A" , x"F" ),
( x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"A" , x"F" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"A" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_5G : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"F" , x"F" , x"3" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"7" , x"7" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"7" , x"7" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"5" , x"5" , x"7" ),
( x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"3" , x"5" , x"0" ),
( x"3" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"0" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"A" , x"A" , x"A" , x"A" , x"A" , x"A" , x"0" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_5B : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"F" , x"F" , x"4" , x"F" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"1" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"4" , x"1" , x"0" ),
( x"4" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_4R : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"F" , x"F" , x"2" , x"F" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"A" , x"A" , x"A" , x"F" , x"F" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"F" , x"F" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"A" , x"A" , x"F" ),
( x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"1" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"B" , x"B" , x"B" , x"B" , x"B" , x"B" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_4G : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"F" , x"F" , x"3" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"7" , x"7" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"7" , x"7" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"5" , x"5" , x"7" ),
( x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"0" ),
( x"3" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_4B : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"F" , x"F" , x"4" , x"F" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"1" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"0" ),
( x"4" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_3R : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"F" , x"F" , x"2" , x"F" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"A" , x"A" , x"A" , x"F" , x"F" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"F" , x"F" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"A" , x"A" , x"F" ),
( x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_3G : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"F" , x"F" , x"3" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"7" , x"7" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"7" , x"7" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"5" , x"5" , x"7" ),
( x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"0" ),
( x"3" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_3B : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"F" , x"F" , x"4" , x"F" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"1" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"0" ),
( x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_2R : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"F" , x"F" , x"2" , x"F" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"A" , x"A" , x"A" , x"F" , x"F" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"F" , x"F" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"A" , x"A" , x"F" ),
( x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_2G : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"F" , x"F" , x"3" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"7" , x"7" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"7" , x"7" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"5" , x"5" , x"7" ),
( x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"0" ),
( x"3" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"0" , x"C" , x"C" , x"C" , x"C" , x"0" , x"C" , x"C" , x"C" , x"C" , x"C" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_2B : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"F" , x"F" , x"4" , x"F" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"1" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"0" ),
( x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_1R : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"F" , x"F" , x"2" , x"F" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"A" , x"A" , x"A" , x"F" , x"F" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"F" , x"2" , x"F" , x"2" , x"F" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"A" , x"F" , x"F" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"A" , x"A" , x"F" ),
( x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"F" ),
( x"2" , x"2" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"A" , x"F" ),
( x"1" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"A" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"1" , x"1" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"E" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"1" , x"2" , x"1" , x"0" , x"0" , x"E" , x"E" , x"E" , x"E" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_1G : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"F" , x"F" , x"3" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"5" , x"7" , x"7" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"F" , x"3" , x"F" , x"3" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"5" , x"7" , x"7" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"5" , x"5" , x"7" ),
( x"0" , x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"7" ),
( x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"0" ),
( x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" ),
( x"2" , x"3" , x"2" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT health_point_1B : ImageMatrix(0 TO 19, 0 TO 43) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"F" , x"F" , x"4" , x"F" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"F" , x"4" , x"F" , x"4" , x"F" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"1" , x"1" , x"2" ),
( x"0" , x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"5" , x"4" , x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"1" , x"2" ),
( x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"1" , x"0" ),
( x"4" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" ),
( x"3" , x"4" , x"3" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"4" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT startR : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"7" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"9" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"9" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"A" , x"6" , x"6" , x"6" , x"2" , x"6" , x"6" , x"6" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"7" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"A" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"6" , x"6" , x"6" , x"6" , x"6" , x"1" , x"6" , x"6" , x"6" , x"6" , x"2" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"4" , x"4" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"9" , x"6" , x"6" , x"6" , x"4" , x"3" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"6" , x"6" , x"6" , x"1" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"6" , x"1" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"0" , x"4" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"E" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"0" , x"1" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"0" , x"1" , x"3" , x"4" , x"4" , x"3" , x"4" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"2" , x"3" , x"4" , x"4" , x"2" , x"0" , x"0" , x"2" , x"3" , x"0" , x"0" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"E" , x"F" , x"F" , x"F" , x"F" , x"9" , x"0" , x"0" , x"B" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"5" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"9" , x"F" , x"F" , x"F" , x"F" , x"F" , x"1" , x"0" , x"0" , x"C" , x"F" , x"A" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"7" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"F" , x"F" , x"E" , x"C" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"8" , x"0" , x"E" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"4" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"1" , x"0" , x"B" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"4" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"A" , x"0" , x"0" , x"0" , x"0" , x"4" , x"F" , x"F" , x"F" , x"F" , x"F" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"8" , x"D" , x"F" , x"F" , x"F" , x"0" , x"0" , x"E" , x"F" , x"F" , x"F" , x"C" , x"C" , x"E" , x"F" , x"E" , x"0" , x"4" , x"6" , x"5" , x"E" , x"F" , x"F" , x"5" , x"6" , x"5" , x"0" , x"6" , x"F" , x"F" , x"6" , x"6" , x"6" , x"6" , x"5" , x"0" , x"4" , x"F" , x"F" , x"7" , x"6" , x"5" , x"9" , x"F" , x"F" , x"2" , x"0" , x"F" , x"F" , x"F" , x"C" , x"C" , x"D" , x"F" , x"F" , x"4" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"7" , x"5" , x"E" , x"F" , x"F" , x"8" , x"0" , x"0" , x"0" , x"7" , x"F" , x"F" , x"8" , x"E" , x"F" , x"A" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"2" , x"0" , x"4" , x"F" , x"F" , x"8" , x"0" , x"C" , x"F" , x"F" , x"0" , x"0" , x"0" , x"B" , x"C" , x"C" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"1" , x"0" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"E" , x"0" , x"0" , x"2" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"5" , x"F" , x"E" , x"0" , x"5" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"4" , x"F" , x"F" , x"D" , x"D" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"A" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"8" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"3" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"1" , x"D" , x"F" , x"F" , x"F" , x"E" , x"5" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"6" , x"0" , x"0" , x"4" , x"F" , x"F" , x"7" , x"5" , x"5" , x"9" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"A" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"8" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"E" , x"E" , x"E" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"4" , x"E" , x"E" , x"F" , x"F" , x"9" , x"1" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"0" , x"4" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"0" , x"F" , x"F" , x"A" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"1" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"8" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"5" , x"F" , x"F" , x"F" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"D" , x"F" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"7" , x"6" , x"7" , x"3" , x"0" , x"0" , x"5" , x"F" , x"F" , x"E" , x"E" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"A" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"1" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"8" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"E" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"E" , x"E" , x"E" , x"F" , x"F" , x"D" , x"0" , x"1" , x"3" , x"2" , x"0" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"8" , x"F" , x"F" , x"3" , x"0" , x"0" , x"F" , x"F" , x"A" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"8" , x"F" , x"E" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"E" , x"1" , x"0" , x"3" , x"F" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"1" , x"F" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"E" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"2" , x"0" , x"3" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"F" , x"E" , x"D" , x"F" , x"F" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"0" , x"C" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"E" , x"F" , x"F" , x"F" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"E" , x"8" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"E" , x"0" , x"1" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"A" , x"1" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"0" , x"5" , x"F" , x"F" , x"2" , x"0" , x"4" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"6" , x"1" , x"0" , x"F" , x"F" , x"E" , x"0" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"1" , x"0" , x"0" , x"0" , x"0" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"A" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"B" , x"C" , x"C" , x"C" , x"C" , x"5" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"6" , x"4" , x"0" , x"0" , x"0" , x"0" , x"3" , x"6" , x"5" , x"5" , x"5" , x"5" , x"5" , x"4" , x"0" , x"2" , x"5" , x"5" , x"1" , x"0" , x"0" , x"2" , x"6" , x"5" , x"0" , x"0" , x"0" , x"4" , x"6" , x"5" , x"5" , x"5" , x"5" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"2" , x"6" , x"5" , x"5" , x"5" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"A" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"3" , x"1" , x"F" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"1" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"1" , x"0" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"1" , x"1" , x"F" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"3" , x"3" , x"F" , x"1" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"1" , x"F" , x"F" , x"1" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"1" , x"2" , x"F" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"3" , x"0" , x"F" , x"F" , x"F" , x"1" , x"1" , x"F" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"1" , x"F" , x"F" , x"F" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"1" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"1" , x"0" , x"0" , x"F" , x"1" , x"1" , x"F" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT startG : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"7" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"9" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"4" , x"1" , x"1" , x"1" , x"0" , x"0" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"8" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"9" , x"6" , x"6" , x"6" , x"2" , x"6" , x"6" , x"6" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"8" , x"2" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"7" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"6" , x"6" , x"6" , x"6" , x"6" , x"1" , x"6" , x"6" , x"6" , x"6" , x"2" , x"3" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"2" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"4" , x"4" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"8" , x"6" , x"6" , x"6" , x"4" , x"3" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"6" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"6" , x"6" , x"6" , x"6" , x"6" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"6" , x"6" , x"6" , x"6" , x"0" , x"0" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"6" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"3" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"3" , x"3" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"3" , x"2" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"2" , x"2" , x"2" , x"3" , x"2" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"4" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"E" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"0" , x"1" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"3" , x"4" , x"4" , x"3" , x"4" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"2" , x"3" , x"4" , x"4" , x"2" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"E" , x"F" , x"F" , x"F" , x"F" , x"8" , x"0" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"5" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"0" , x"0" , x"0" , x"9" , x"F" , x"F" , x"F" , x"F" , x"E" , x"1" , x"1" , x"1" , x"B" , x"F" , x"9" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"7" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"4" , x"F" , x"F" , x"E" , x"C" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"7" , x"0" , x"E" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"4" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"1" , x"0" , x"A" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"4" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"0" , x"1" , x"1" , x"0" , x"4" , x"E" , x"F" , x"F" , x"F" , x"F" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"E" , x"F" , x"7" , x"D" , x"F" , x"F" , x"F" , x"0" , x"0" , x"E" , x"F" , x"F" , x"F" , x"C" , x"C" , x"E" , x"F" , x"D" , x"0" , x"4" , x"6" , x"5" , x"E" , x"F" , x"E" , x"5" , x"6" , x"5" , x"0" , x"6" , x"F" , x"F" , x"6" , x"6" , x"6" , x"6" , x"5" , x"0" , x"4" , x"F" , x"F" , x"7" , x"6" , x"5" , x"8" , x"F" , x"F" , x"2" , x"0" , x"F" , x"F" , x"F" , x"C" , x"C" , x"D" , x"F" , x"F" , x"4" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"7" , x"5" , x"E" , x"F" , x"F" , x"7" , x"0" , x"0" , x"0" , x"7" , x"F" , x"F" , x"7" , x"D" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"E" , x"2" , x"0" , x"4" , x"F" , x"F" , x"7" , x"0" , x"C" , x"F" , x"F" , x"0" , x"0" , x"0" , x"B" , x"C" , x"C" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"1" , x"0" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"E" , x"F" , x"D" , x"0" , x"0" , x"2" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"0" , x"0" , x"5" , x"F" , x"E" , x"0" , x"5" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"4" , x"F" , x"F" , x"D" , x"D" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"F" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"0" , x"4" , x"F" , x"F" , x"1" , x"0" , x"E" , x"F" , x"9" , x"0" , x"1" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"7" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"3" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"1" , x"D" , x"F" , x"F" , x"F" , x"E" , x"5" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"1" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"6" , x"0" , x"0" , x"4" , x"F" , x"F" , x"7" , x"5" , x"5" , x"9" , x"F" , x"F" , x"1" , x"0" , x"E" , x"F" , x"9" , x"0" , x"1" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"E" , x"E" , x"E" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"4" , x"E" , x"E" , x"F" , x"F" , x"9" , x"1" , x"0" , x"0" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"0" , x"4" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"1" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"1" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"5" , x"F" , x"F" , x"E" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"D" , x"F" , x"F" , x"8" , x"0" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"1" , x"6" , x"F" , x"F" , x"7" , x"6" , x"7" , x"3" , x"0" , x"1" , x"5" , x"E" , x"F" , x"E" , x"E" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"1" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"E" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"E" , x"E" , x"E" , x"F" , x"F" , x"D" , x"0" , x"1" , x"3" , x"2" , x"0" , x"0" , x"0" , x"D" , x"F" , x"8" , x"0" , x"0" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"4" , x"F" , x"F" , x"2" , x"0" , x"7" , x"F" , x"F" , x"3" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"0" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"C" , x"1" , x"0" , x"3" , x"E" , x"F" , x"8" , x"0" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"F" , x"1" , x"1" , x"2" , x"2" , x"2" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"1" , x"F" , x"F" , x"E" , x"1" , x"0" , x"E" , x"F" , x"E" , x"0" , x"1" , x"4" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"2" , x"0" , x"3" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"F" , x"C" , x"C" , x"F" , x"F" , x"F" , x"9" , x"0" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"C" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"0" , x"C" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"D" , x"F" , x"F" , x"F" , x"F" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"E" , x"E" , x"C" , x"7" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"1" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"1" , x"0" , x"0" , x"1" , x"0" , x"E" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"0" , x"4" , x"F" , x"F" , x"2" , x"0" , x"0" , x"5" , x"F" , x"E" , x"2" , x"0" , x"4" , x"B" , x"F" , x"F" , x"F" , x"F" , x"F" , x"6" , x"1" , x"0" , x"E" , x"F" , x"D" , x"0" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"1" , x"0" , x"0" , x"0" , x"0" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"B" , x"C" , x"C" , x"C" , x"C" , x"5" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"3" , x"6" , x"4" , x"0" , x"0" , x"1" , x"0" , x"3" , x"6" , x"5" , x"5" , x"5" , x"5" , x"5" , x"4" , x"0" , x"2" , x"5" , x"5" , x"1" , x"0" , x"0" , x"2" , x"6" , x"5" , x"0" , x"0" , x"0" , x"4" , x"6" , x"5" , x"5" , x"5" , x"5" , x"0" , x"0" , x"1" , x"4" , x"6" , x"3" , x"0" , x"2" , x"6" , x"5" , x"5" , x"5" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"2" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"1" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"F" , x"F" , x"3" , x"1" , x"F" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"1" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"1" , x"0" , x"F" , x"F" , x"F" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"1" , x"1" , x"F" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"3" , x"3" , x"F" , x"1" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"1" , x"F" , x"F" , x"1" , x"0" , x"0" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"1" , x"2" , x"F" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"3" , x"0" , x"F" , x"F" , x"F" , x"1" , x"1" , x"F" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"0" , x"2" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"1" , x"F" , x"F" , x"F" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"1" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"2" , x"1" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"1" , x"0" , x"0" , x"F" , x"1" , x"1" , x"F" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"3" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"1" , x"2" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"2" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"4" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);

CONSTANT startB : ImageMatrix(0 TO 74, 0 TO 99) := (
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"3" , x"1" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"0" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"3" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"1" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"2" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"4" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"1" , x"1" , x"2" , x"1" , x"3" , x"3" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"2" , x"3" , x"5" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"3" , x"2" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"4" , x"7" , x"7" , x"7" , x"7" , x"7" , x"4" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"2" , x"2" , x"2" , x"3" , x"2" , x"1" , x"2" , x"2" , x"2" , x"3" , x"5" , x"3" , x"4" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"4" , x"4" , x"1" , x"2" , x"1" , x"0" , x"1" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"4" , x"6" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"4" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"4" , x"2" , x"4" , x"6" , x"4" , x"4" , x"5" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"4" , x"2" , x"2" , x"0" , x"1" , x"0" , x"2" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"6" , x"7" , x"7" , x"7" , x"7" , x"6" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"2" , x"3" , x"2" , x"3" , x"1" , x"2" , x"3" , x"3" , x"3" , x"5" , x"6" , x"5" , x"6" , x"4" , x"3" , x"4" , x"4" , x"3" , x"3" , x"4" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"7" , x"7" , x"7" , x"8" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"2" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"4" , x"5" , x"3" , x"3" , x"3" , x"2" , x"1" , x"5" , x"4" , x"3" , x"4" , x"3" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"1" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"0" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"9" , x"7" , x"7" , x"7" , x"4" , x"7" , x"7" , x"7" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"2" , x"3" , x"3" , x"4" , x"3" , x"4" , x"7" , x"4" , x"3" , x"3" , x"4" , x"3" , x"4" , x"5" , x"6" , x"2" , x"3" , x"4" , x"3" , x"4" , x"3" , x"1" , x"4" , x"0" , x"0" , x"1" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"7" , x"7" , x"7" , x"7" , x"7" , x"2" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"1" , x"7" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"9" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"3" , x"4" , x"4" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"2" , x"5" , x"6" , x"6" , x"6" , x"6" , x"4" , x"4" , x"2" , x"3" , x"2" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"1" , x"3" , x"3" , x"2" , x"2" , x"3" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"7" , x"7" , x"7" , x"7" , x"6" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"1" , x"2" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"5" , x"6" , x"6" , x"6" , x"2" , x"1" , x"3" , x"4" , x"1" , x"2" , x"1" , x"2" , x"0" , x"1" , x"0" , x"0" , x"2" , x"2" , x"1" , x"3" , x"4" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"0" , x"1" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"2" , x"7" , x"7" , x"7" , x"7" , x"7" , x"3" , x"7" , x"7" , x"7" , x"7" , x"4" , x"4" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"2" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"4" , x"5" , x"6" , x"6" , x"4" , x"1" , x"4" , x"3" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"3" , x"4" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"3" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"4" , x"5" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"6" , x"5" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"1" , x"1" , x"3" , x"3" , x"2" , x"2" , x"1" , x"2" , x"4" , x"2" , x"3" , x"1" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"5" , x"4" , x"3" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"1" , x"3" , x"1" , x"3" , x"3" , x"2" , x"3" , x"4" , x"2" , x"2" , x"3" , x"3" , x"5" , x"6" , x"6" , x"4" , x"3" , x"3" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"4" , x"2" , x"3" , x"5" , x"4" , x"3" , x"3" , x"2" , x"1" , x"0" , x"1" , x"0" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"7" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"3" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"5" , x"6" , x"6" , x"6" , x"4" , x"2" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"5" , x"4" , x"4" , x"3" , x"3" , x"2" , x"2" , x"1" , x"0" , x"1" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"7" , x"7" , x"7" , x"7" , x"7" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"0" , x"2" , x"0" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"4" , x"1" , x"2" , x"4" , x"5" , x"6" , x"6" , x"6" , x"4" , x"3" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"5" , x"4" , x"2" , x"3" , x"1" , x"1" , x"2" , x"3" , x"1" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"7" , x"7" , x"7" , x"0" , x"0" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"1" , x"3" , x"4" , x"3" , x"5" , x"6" , x"6" , x"4" , x"4" , x"5" , x"2" , x"1" , x"0" , x"0" , x"2" , x"2" , x"2" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"5" , x"3" , x"4" , x"4" , x"4" , x"2" , x"2" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" ),
( x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"4" , x"7" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"3" , x"2" , x"1" , x"3" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"5" , x"6" , x"5" , x"5" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"4" , x"2" , x"2" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"3" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"5" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"3" , x"2" , x"2" , x"2" , x"2" , x"3" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"2" , x"2" , x"1" , x"1" , x"2" , x"2" , x"3" , x"4" , x"4" , x"3" , x"4" , x"5" , x"5" , x"4" , x"2" , x"3" , x"2" , x"1" , x"1" , x"3" , x"3" , x"1" , x"0" , x"0" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"7" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"3" , x"1" , x"3" , x"2" , x"3" , x"2" , x"2" , x"1" , x"1" , x"1" , x"3" , x"3" , x"2" , x"3" , x"3" , x"1" , x"0" , x"2" , x"1" , x"1" , x"2" , x"2" , x"2" , x"4" , x"4" , x"4" , x"4" , x"3" , x"5" , x"4" , x"3" , x"3" , x"2" , x"3" , x"1" , x"2" , x"3" , x"1" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"3" , x"2" , x"3" , x"2" , x"3" , x"4" , x"1" , x"0" , x"0" , x"0" , x"2" , x"3" , x"2" , x"3" , x"4" , x"3" , x"4" , x"4" , x"3" , x"4" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"3" , x"2" , x"0" , x"2" , x"2" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"5" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"3" , x"3" , x"2" , x"3" , x"4" , x"0" , x"0" , x"1" , x"3" , x"3" , x"3" , x"3" , x"3" , x"5" , x"4" , x"4" , x"3" , x"3" , x"0" , x"0" , x"2" , x"2" , x"3" , x"3" , x"4" , x"3" , x"4" , x"4" , x"3" , x"2" , x"1" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"3" , x"2" , x"2" , x"3" , x"3" , x"2" , x"1" , x"1" , x"2" , x"1" , x"2" , x"3" , x"3" , x"1" , x"3" , x"6" , x"5" , x"4" , x"3" , x"2" , x"0" , x"0" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"1" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"0" , x"0" , x"0" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"2" , x"3" , x"3" , x"2" , x"1" , x"0" , x"1" , x"2" , x"0" , x"3" , x"4" , x"3" , x"3" , x"4" , x"4" , x"5" , x"4" , x"2" , x"1" , x"0" , x"0" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"2" , x"3" , x"4" , x"4" , x"1" , x"3" , x"3" , x"1" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"1" , x"3" , x"3" , x"0" , x"1" , x"2" , x"3" , x"2" , x"1" , x"4" , x"4" , x"4" , x"6" , x"5" , x"2" , x"4" , x"3" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"3" , x"4" , x"4" , x"3" , x"4" , x"4" , x"3" , x"4" , x"1" , x"1" , x"3" , x"2" , x"1" , x"2" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"1" , x"2" , x"2" , x"3" , x"4" , x"4" , x"3" , x"3" , x"4" , x"3" , x"5" , x"3" , x"1" , x"2" , x"1" , x"4" , x"2" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"2" , x"1" , x"0" , x"0" , x"2" , x"3" , x"1" , x"3" , x"3" , x"3" , x"4" , x"3" , x"1" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"2" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"E" , x"F" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"4" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"4" , x"4" , x"4" , x"4" , x"2" , x"0" , x"2" , x"3" , x"4" , x"4" , x"4" , x"2" , x"2" , x"2" , x"2" , x"3" , x"4" , x"5" , x"4" , x"4" , x"4" , x"4" , x"4" , x"2" , x"0" , x"0" , x"0" , x"2" , x"4" , x"4" , x"4" , x"4" , x"5" , x"4" , x"2" , x"3" , x"4" , x"4" , x"5" , x"3" , x"4" , x"4" , x"4" , x"4" , x"2" , x"2" , x"0" , x"1" , x"2" , x"1" , x"0" , x"1" , x"2" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"1" , x"E" , x"F" , x"E" , x"E" , x"F" , x"7" , x"1" , x"0" , x"9" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"E" , x"A" , x"1" , x"7" , x"C" , x"E" , x"E" , x"E" , x"E" , x"E" , x"A" , x"1" , x"5" , x"C" , x"E" , x"E" , x"E" , x"E" , x"E" , x"A" , x"0" , x"0" , x"0" , x"0" , x"8" , x"C" , x"E" , x"E" , x"E" , x"B" , x"2" , x"2" , x"2" , x"A" , x"F" , x"9" , x"1" , x"6" , x"C" , x"E" , x"E" , x"E" , x"E" , x"6" , x"0" , x"1" , x"0" , x"0" , x"2" , x"1" , x"4" , x"E" , x"F" , x"E" , x"C" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"F" , x"F" , x"E" , x"F" , x"E" , x"0" , x"0" , x"C" , x"E" , x"F" , x"F" , x"F" , x"F" , x"E" , x"E" , x"7" , x"0" , x"E" , x"F" , x"F" , x"E" , x"F" , x"F" , x"E" , x"F" , x"E" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"5" , x"F" , x"E" , x"F" , x"F" , x"F" , x"E" , x"E" , x"A" , x"2" , x"0" , x"9" , x"E" , x"E" , x"F" , x"F" , x"F" , x"E" , x"A" , x"4" , x"2" , x"E" , x"F" , x"D" , x"0" , x"7" , x"F" , x"E" , x"F" , x"F" , x"F" , x"F" , x"9" , x"0" , x"2" , x"2" , x"1" , x"4" , x"E" , x"F" , x"F" , x"F" , x"F" , x"5" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"D" , x"F" , x"7" , x"D" , x"F" , x"F" , x"F" , x"0" , x"0" , x"E" , x"F" , x"F" , x"F" , x"C" , x"C" , x"D" , x"F" , x"D" , x"0" , x"5" , x"6" , x"5" , x"E" , x"F" , x"E" , x"5" , x"6" , x"5" , x"0" , x"6" , x"F" , x"E" , x"6" , x"6" , x"6" , x"6" , x"5" , x"0" , x"5" , x"F" , x"E" , x"6" , x"6" , x"5" , x"7" , x"E" , x"E" , x"2" , x"1" , x"E" , x"F" , x"F" , x"C" , x"C" , x"D" , x"E" , x"F" , x"4" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"6" , x"5" , x"E" , x"F" , x"E" , x"7" , x"0" , x"1" , x"1" , x"6" , x"F" , x"F" , x"7" , x"D" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"B" , x"2" , x"0" , x"4" , x"F" , x"F" , x"7" , x"0" , x"C" , x"F" , x"E" , x"0" , x"0" , x"0" , x"B" , x"C" , x"C" , x"0" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"E" , x"2" , x"0" , x"0" , x"4" , x"F" , x"E" , x"2" , x"1" , x"E" , x"F" , x"D" , x"0" , x"0" , x"2" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"D" , x"F" , x"E" , x"0" , x"1" , x"1" , x"5" , x"E" , x"E" , x"0" , x"5" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"4" , x"F" , x"E" , x"D" , x"D" , x"3" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"3" , x"3" , x"1" , x"7" , x"F" , x"E" , x"1" , x"4" , x"4" , x"4" , x"3" , x"1" , x"5" , x"F" , x"E" , x"2" , x"0" , x"1" , x"5" , x"F" , x"E" , x"2" , x"0" , x"E" , x"F" , x"9" , x"0" , x"3" , x"5" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"2" , x"0" , x"0" , x"7" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"6" , x"F" , x"D" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"3" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"2" , x"D" , x"F" , x"F" , x"F" , x"D" , x"5" , x"3" , x"0" , x"0" , x"1" , x"1" , x"0" , x"D" , x"F" , x"E" , x"0" , x"2" , x"4" , x"2" , x"7" , x"F" , x"F" , x"F" , x"F" , x"E" , x"6" , x"1" , x"1" , x"5" , x"F" , x"E" , x"6" , x"5" , x"5" , x"8" , x"E" , x"E" , x"2" , x"0" , x"E" , x"F" , x"9" , x"0" , x"3" , x"4" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"E" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"F" , x"F" , x"F" , x"E" , x"E" , x"E" , x"E" , x"F" , x"D" , x"0" , x"0" , x"1" , x"4" , x"E" , x"E" , x"F" , x"F" , x"8" , x"1" , x"0" , x"0" , x"2" , x"1" , x"D" , x"F" , x"E" , x"0" , x"3" , x"4" , x"2" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"1" , x"2" , x"5" , x"F" , x"E" , x"F" , x"F" , x"F" , x"F" , x"E" , x"C" , x"0" , x"1" , x"E" , x"F" , x"9" , x"0" , x"2" , x"5" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"1" , x"6" , x"F" , x"E" , x"2" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"1" , x"0" , x"0" , x"1" , x"5" , x"E" , x"F" , x"E" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"B" , x"D" , x"E" , x"F" , x"7" , x"0" , x"2" , x"3" , x"1" , x"D" , x"F" , x"E" , x"0" , x"2" , x"3" , x"3" , x"7" , x"F" , x"E" , x"6" , x"6" , x"6" , x"3" , x"1" , x"3" , x"5" , x"C" , x"E" , x"E" , x"E" , x"E" , x"F" , x"F" , x"0" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"2" , x"4" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"1" , x"6" , x"F" , x"E" , x"2" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"5" , x"F" , x"F" , x"D" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"6" , x"5" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"E" , x"E" , x"E" , x"E" , x"F" , x"F" , x"D" , x"0" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"D" , x"F" , x"7" , x"0" , x"2" , x"3" , x"1" , x"D" , x"F" , x"E" , x"0" , x"2" , x"3" , x"2" , x"6" , x"F" , x"E" , x"0" , x"0" , x"0" , x"0" , x"3" , x"3" , x"5" , x"E" , x"E" , x"2" , x"0" , x"7" , x"F" , x"E" , x"3" , x"0" , x"0" , x"E" , x"F" , x"9" , x"0" , x"1" , x"4" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"1" , x"0" , x"0" , x"7" , x"F" , x"E" , x"0" , x"0" , x"0" , x"5" , x"E" , x"F" , x"D" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"5" , x"4" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"A" , x"2" , x"0" , x"3" , x"E" , x"F" , x"7" , x"0" , x"2" , x"2" , x"2" , x"D" , x"F" , x"E" , x"0" , x"2" , x"3" , x"1" , x"6" , x"F" , x"E" , x"2" , x"3" , x"4" , x"4" , x"4" , x"1" , x"5" , x"E" , x"E" , x"2" , x"0" , x"2" , x"E" , x"F" , x"C" , x"2" , x"1" , x"E" , x"F" , x"D" , x"0" , x"2" , x"4" , x"E" , x"E" , x"3" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"2" , x"0" , x"3" , x"E" , x"F" , x"E" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"F" , x"F" , x"D" , x"0" , x"0" , x"0" , x"E" , x"F" , x"D" , x"0" , x"C" , x"F" , x"E" , x"A" , x"A" , x"E" , x"E" , x"F" , x"8" , x"0" , x"2" , x"3" , x"1" , x"D" , x"F" , x"E" , x"0" , x"3" , x"3" , x"1" , x"6" , x"E" , x"F" , x"E" , x"E" , x"E" , x"E" , x"A" , x"1" , x"5" , x"E" , x"E" , x"2" , x"0" , x"0" , x"C" , x"F" , x"E" , x"2" , x"1" , x"E" , x"E" , x"B" , x"E" , x"E" , x"E" , x"E" , x"F" , x"3" , x"0" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"E" , x"E" , x"E" , x"E" , x"F" , x"E" , x"1" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"E" , x"E" , x"A" , x"7" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"F" , x"F" , x"D" , x"0" , x"1" , x"0" , x"E" , x"F" , x"D" , x"0" , x"1" , x"C" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"2" , x"0" , x"0" , x"2" , x"1" , x"D" , x"F" , x"F" , x"0" , x"1" , x"1" , x"1" , x"7" , x"F" , x"F" , x"F" , x"F" , x"F" , x"F" , x"E" , x"0" , x"5" , x"F" , x"F" , x"2" , x"0" , x"0" , x"5" , x"D" , x"C" , x"2" , x"1" , x"4" , x"A" , x"F" , x"F" , x"F" , x"F" , x"F" , x"6" , x"1" , x"1" , x"E" , x"F" , x"D" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"8" , x"1" , x"0" , x"0" , x"0" , x"0" , x"6" , x"F" , x"F" , x"F" , x"F" , x"F" , x"9" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"0" , x"4" , x"6" , x"3" , x"0" , x"0" , x"B" , x"C" , x"C" , x"C" , x"C" , x"5" , x"2" , x"0" , x"0" , x"1" , x"2" , x"1" , x"3" , x"6" , x"4" , x"0" , x"1" , x"3" , x"2" , x"4" , x"6" , x"5" , x"5" , x"5" , x"5" , x"5" , x"5" , x"0" , x"4" , x"5" , x"5" , x"1" , x"0" , x"1" , x"4" , x"6" , x"5" , x"0" , x"2" , x"2" , x"4" , x"6" , x"5" , x"5" , x"5" , x"5" , x"0" , x"0" , x"3" , x"5" , x"6" , x"3" , x"0" , x"2" , x"6" , x"5" , x"5" , x"5" , x"5" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"5" , x"5" , x"5" , x"5" , x"5" , x"3" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"1" , x"0" , x"1" , x"0" , x"1" , x"3" , x"3" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"1" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"1" , x"2" , x"1" , x"0" , x"2" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"4" , x"4" , x"3" , x"4" , x"3" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"3" , x"2" , x"3" , x"4" , x"4" , x"3" , x"1" , x"3" , x"4" , x"5" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"1" , x"2" , x"2" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"2" , x"2" , x"0" , x"1" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"3" , x"3" , x"4" , x"4" , x"5" , x"4" , x"4" , x"3" , x"1" , x"3" , x"4" , x"3" , x"3" , x"3" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"2" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"1" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"5" , x"4" , x"4" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"3" , x"4" , x"3" , x"2" , x"3" , x"4" , x"6" , x"6" , x"5" , x"3" , x"3" , x"3" , x"1" , x"3" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"1" , x"2" , x"2" , x"1" , x"2" , x"1" , x"3" , x"4" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"2" , x"3" , x"2" , x"3" , x"3" , x"4" , x"5" , x"3" , x"3" , x"3" , x"4" , x"4" , x"3" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"2" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"4" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"3" , x"3" , x"4" , x"3" , x"3" , x"3" , x"2" , x"4" , x"4" , x"3" , x"4" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"3" , x"3" , x"5" , x"4" , x"5" , x"4" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"4" , x"3" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"6" , x"6" , x"4" , x"4" , x"2" , x"2" , x"1" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"5" , x"5" , x"4" , x"3" , x"3" , x"2" , x"3" , x"2" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"3" , x"2" , x"3" , x"4" , x"5" , x"6" , x"4" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"2" , x"4" , x"4" , x"4" , x"4" , x"6" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"0" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"2" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"2" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"1" , x"3" , x"5" , x"5" , x"5" , x"3" , x"3" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"2" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"5" , x"5" , x"5" , x"4" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"5" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"0" , x"1" , x"2" , x"3" , x"2" , x"3" , x"2" , x"4" , x"5" , x"3" , x"2" , x"3" , x"2" , x"2" , x"0" , x"1" , x"3" , x"1" , x"0" , x"0" , x"2" , x"3" , x"3" , x"3" , x"4" , x"5" , x"4" , x"4" , x"5" , x"3" , x"3" , x"4" , x"2" , x"1" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"1" , x"3" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"2" , x"2" , x"4" , x"5" , x"4" , x"0" , x"1" , x"2" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"5" , x"4" , x"2" , x"3" , x"1" , x"1" , x"2" , x"3" , x"1" , x"2" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"3" , x"3" , x"2" , x"3" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"0" , x"1" , x"2" , x"1" , x"2" , x"3" , x"2" , x"1" , x"2" , x"2" , x"4" , x"4" , x"4" , x"3" , x"3" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"2" , x"1" , x"0" , x"1" , x"2" , x"2" , x"3" , x"4" , x"4" , x"5" , x"4" , x"5" , x"4" , x"3" , x"3" , x"3" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"3" , x"3" , x"2" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"2" , x"1" , x"2" , x"1" , x"1" , x"2" , x"1" , x"2" , x"3" , x"3" , x"4" , x"5" , x"5" , x"4" , x"2" , x"2" , x"1" , x"1" , x"0" , x"2" , x"1" , x"2" , x"1" , x"1" , x"2" , x"2" , x"1" , x"3" , x"4" , x"4" , x"4" , x"4" , x"5" , x"3" , x"2" , x"3" , x"3" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"2" , x"3" , x"3" , x"1" , x"2" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"3" , x"3" , x"4" , x"3" , x"4" , x"5" , x"4" , x"3" , x"3" , x"1" , x"1" , x"2" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"1" , x"3" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"2" , x"3" , x"2" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"3" , x"2" , x"2" , x"3" , x"3" , x"2" , x"3" , x"4" , x"4" , x"3" , x"2" , x"3" , x"3" , x"1" , x"1" , x"2" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"5" , x"9" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"5" , x"3" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"3" , x"3" , x"3" , x"4" , x"3" , x"3" , x"4" , x"3" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"2" , x"3" , x"5" , x"5" , x"4" , x"4" , x"3" , x"1" , x"1" , x"0" , x"F" , x"F" , x"3" , x"3" , x"F" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"F" , x"1" , x"1" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"1" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"1" , x"0" , x"F" , x"F" , x"F" , x"3" , x"3" , x"3" , x"3" , x"3" , x"4" , x"5" , x"3" , x"3" , x"4" , x"1" , x"2" , x"3" , x"1" , x"1" , x"1" , x"2" , x"1" , x"1" , x"2" , x"3" , x"3" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"3" , x"3" , x"3" , x"2" , x"3" , x"3" , x"5" , x"5" , x"5" , x"3" , x"2" , x"2" , x"0" , x"0" , x"F" , x"2" , x"F" , x"1" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"0" , x"0" , x"1" , x"0" , x"F" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"1" , x"F" , x"1" , x"1" , x"F" , x"0" , x"F" , x"2" , x"F" , x"0" , x"F" , x"0" , x"0" , x"3" , x"3" , x"3" , x"4" , x"5" , x"5" , x"4" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"2" , x"1" , x"3" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"2" , x"3" , x"3" , x"3" , x"3" , x"4" , x"3" , x"4" , x"6" , x"5" , x"4" , x"2" , x"2" , x"1" , x"0" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"3" , x"3" , x"F" , x"1" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"1" , x"1" , x"F" , x"F" , x"1" , x"0" , x"1" , x"0" , x"F" , x"F" , x"F" , x"0" , x"F" , x"1" , x"F" , x"0" , x"F" , x"1" , x"1" , x"F" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"F" , x"0" , x"4" , x"4" , x"5" , x"5" , x"5" , x"5" , x"3" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"3" , x"3" , x"1" , x"2" , x"3" , x"4" , x"4" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"F" , x"F" , x"3" , x"1" , x"F" , x"F" , x"F" , x"1" , x"1" , x"F" , x"1" , x"2" , x"0" , x"1" , x"F" , x"F" , x"1" , x"0" , x"F" , x"F" , x"1" , x"0" , x"0" , x"0" , x"0" , x"F" , x"0" , x"F" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"F" , x"0" , x"0" , x"4" , x"4" , x"5" , x"4" , x"4" , x"2" , x"1" , x"2" , x"4" , x"4" , x"3" , x"4" , x"2" , x"3" , x"3" , x"1" , x"0" , x"1" , x"0" , x"1" , x"3" , x"2" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"2" , x"3" , x"3" , x"3" , x"5" , x"5" , x"5" , x"5" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"F" , x"1" , x"1" , x"1" , x"F" , x"0" , x"1" , x"F" , x"1" , x"F" , x"F" , x"F" , x"1" , x"F" , x"F" , x"1" , x"F" , x"F" , x"F" , x"1" , x"0" , x"0" , x"F" , x"F" , x"F" , x"1" , x"0" , x"F" , x"0" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"0" , x"0" , x"F" , x"F" , x"F" , x"4" , x"5" , x"4" , x"4" , x"2" , x"1" , x"1" , x"3" , x"5" , x"3" , x"4" , x"4" , x"3" , x"5" , x"4" , x"2" , x"3" , x"1" , x"0" , x"0" , x"1" , x"3" , x"3" , x"1" , x"0" , x"2" , x"2" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"2" , x"3" , x"3" , x"4" , x"5" , x"4" , x"4" , x"4" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"0" , x"0" , x"1" , x"F" , x"3" , x"2" , x"2" , x"F" , x"3" , x"3" , x"F" , x"3" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"3" , x"5" , x"5" , x"2" , x"1" , x"2" , x"3" , x"3" , x"4" , x"5" , x"4" , x"4" , x"4" , x"4" , x"6" , x"4" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"2" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"2" , x"2" , x"3" , x"2" , x"4" , x"6" , x"5" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"1" , x"0" , x"1" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"3" , x"3" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"1" , x"1" , x"1" , x"1" , x"3" , x"4" , x"4" , x"3" , x"2" , x"1" , x"2" , x"4" , x"5" , x"4" , x"4" , x"4" , x"5" , x"4" , x"2" , x"4" , x"5" , x"4" , x"2" , x"1" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"2" , x"2" , x"2" , x"4" , x"5" , x"6" , x"3" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"1" , x"2" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"3" , x"4" , x"4" , x"3" , x"3" , x"1" , x"1" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"0" , x"1" , x"2" , x"3" , x"4" , x"5" , x"4" , x"3" , x"1" , x"1" , x"2" , x"4" , x"4" , x"3" , x"0" , x"1" , x"2" , x"2" , x"3" , x"3" , x"4" , x"4" , x"3" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"3" , x"2" , x"5" , x"5" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"0" , x"1" , x"3" , x"3" , x"4" , x"4" , x"4" , x"2" , x"1" , x"2" , x"3" , x"3" , x"2" , x"0" , x"0" , x"0" , x"2" , x"1" , x"3" , x"5" , x"3" , x"4" , x"3" , x"2" , x"1" , x"0" , x"2" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"2" , x"3" , x"3" , x"4" , x"3" , x"3" , x"3" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"2" , x"3" , x"4" , x"4" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"0" , x"2" , x"1" , x"2" , x"1" , x"3" , x"4" , x"4" , x"3" , x"4" , x"2" , x"2" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"3" , x"3" , x"3" , x"3" , x"3" , x"3" , x"2" , x"3" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"3" , x"1" , x"1" , x"2" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"2" , x"3" , x"1" , x"1" , x"0" , x"3" , x"1" , x"0" , x"1" , x"4" , x"3" , x"3" , x"4" , x"1" , x"0" , x"0" , x"0" , x"1" , x"3" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"3" , x"2" , x"0" , x"1" , x"3" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"1" , x"0" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"2" , x"4" , x"3" , x"3" , x"3" , x"2" , x"3" , x"2" , x"2" , x"2" , x"3" , x"2" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"3" , x"1" , x"0" , x"2" , x"0" , x"1" , x"1" , x"0" , x"1" , x"3" , x"4" , x"3" , x"3" , x"2" , x"2" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"2" , x"1" , x"2" , x"3" , x"5" , x"4" , x"4" , x"4" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"2" , x"1" , x"3" , x"3" , x"2" , x"1" , x"0" , x"2" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"2" , x"4" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"2" , x"3" , x"2" , x"2" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"1" , x"2" , x"3" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"1" , x"1" , x"2" , x"0" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"2" , x"2" , x"2" , x"1" , x"0" , x"1" , x"1" , x"0" , x"0" , x"2" , x"1" , x"2" , x"3" , x"3" , x"2" , x"0" , x"1" , x"3" , x"4" , x"3" , x"2" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"1" , x"1" , x"0" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"2" , x"0" , x"0" , x"1" , x"1" , x"2" , x"2" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"4" , x"4" , x"4" , x"1" , x"1" , x"2" , x"2" , x"2" , x"2" , x"3" , x"3" , x"3" , x"4" , x"3" , x"1" , x"0" , x"2" , x"2" , x"3" , x"4" , x"1" , x"1" , x"3" , x"1" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"1" , x"1" , x"1" , x"0" , x"2" , x"0" , x"1" , x"2" , x"1" , x"2" , x"2" , x"3" , x"3" , x"4" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"1" , x"2" , x"2" , x"0" , x"0" , x"1" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"4" , x"3" , x"3" , x"3" , x"4" , x"1" , x"2" , x"1" , x"0" , x"0" , x"2" , x"3" , x"3" , x"1" , x"0" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"2" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"1" , x"4" , x"3" , x"2" , x"2" , x"3" , x"3" , x"2" , x"2" , x"3" , x"1" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"1" , x"1" , x"3" , x"3" , x"4" , x"4" , x"3" , x"4" , x"4" , x"4" , x"4" , x"3" , x"4" , x"4" , x"3" , x"2" , x"1" , x"1" , x"0" , x"0" , x"0" , x"3" , x"2" , x"2" , x"2" , x"0" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"2" , x"2" , x"2" , x"4" , x"3" , x"2" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"1" , x"2" , x"2" , x"2" , x"3" , x"4" , x"4" , x"4" , x"4" , x"4" , x"4" , x"3" , x"3" , x"3" , x"2" , x"1" , x"0" , x"0" , x"0" , x"0" , x"1" , x"4" , x"2" , x"2" , x"2" , x"3" , x"1" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" ),
( x"0" , x"0" , x"0" , x"0" , x"1" , x"2" , x"3" , x"2" , x"2" , x"3" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"2" , x"3" , x"1" , x"0" , x"2" , x"0" , x"1" , x"0" , x"0" , x"1" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"1" , x"1" , x"0" , x"1" , x"1" , x"2" , x"2" , x"3" , x"3" , x"3" , x"3" , x"2" , x"2" , x"2" , x"2" , x"1" , x"2" , x"0" , x"0" , x"0" , x"1" , x"3" , x"4" , x"3" , x"1" , x"1" , x"2" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" , x"0" )
);


END ImagePackage;